
module top;
    `include "foo.svh"
endmodule
